module alu_TB();
reg in_TB,
 wire ou_TB


//internal_signals
  reg name_TB;

alu alu_inst(
.in(in_TB),
.ou(ou_TB)
);

endmodule
