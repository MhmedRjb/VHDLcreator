module alu(
  input wire a,
  input wire B,
  input wire C,
  input wire D,
  output reg OB,
  output reg hgf,
  output reg gf
);

//internal_signals
  wire fsdgsyu;

endmodule
