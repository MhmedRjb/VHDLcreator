module alu(
  input wire in,
  output reg ou
);

//internal_signals
  wire name;

endmodule
